module fv_uC_8bits (
    // BlackBox
    input  logic         clk,
    input  logic         clk_valid,
    input  logic         arst_n,
    input  logic [15:0]  flash_data,
    input  logic [7:0]   in,
    input  logic [7:0]   out0, out1,
    input  logic [11:0]  pc_out,

    input  logic         bootstrapping,
    input  logic         cu_state,
    input  logic         equal_flag, carry_flag,
    input  logic         out_select,

    // WhiteBox
    input  logic         equal, carry_out,
    input  logic [7:0]   alu_result,
    input  logic [7:0]   alu_a, alu_b,
    input  logic [2:0]   alu_opcode,

    input  logic         pc_load,
    input  logic [11:0]  pc_next,
    input  logic         pc_inc, 

    input  logic         sram_write_en,
    input  logic [5:0]   sram_addr,
    input  logic [7:0]   sram_data_out,
    input  logic [7:0]   sram_data_in
);
    `include "includes.vh"

    localparam int DELAY = 2;

    `ASM(uC_8bits, clk_valid,
        1'b1 |->, clk_valid ==  1'b1 
    )

    // =============================== ADD assert BlackBox 
    logic [8:0] add_result;
    logic [7:0] add_a, add_b;
    sequence add_sequence;
        (flash_data == {8'h61, add_a}) ##DELAY
        (flash_data == {8'h62, add_b}) ##DELAY
        (flash_data == 16'h8312);// SUM
    endsequence

    logic [7:0] add_a_reg, add_b_reg;
    bus_shift #(.DELAY(5), .WIDTH(8)) add_a_shifting (
        .clk(clk),
        .arst_n(arst_n),
        .in(add_a),
        .out(add_a_reg)
    );
    bus_shift #(.DELAY(3), .WIDTH(8)) add_b_shifting (
        .clk(clk),
        .arst_n(arst_n),
        .in(add_b),
        .out(add_b_reg)
    );

    assign add_result = add_b_reg + add_a_reg;

    property p_exec_sum_from_reset;
    @(posedge clk) disable iff (!arst_n)
        $rose(arst_n) |-> add_sequence |=> (alu_opcode==3'b000 && alu_result==add_result[7:0]);
    endproperty


    // =============================== SUB assert BlackBox 
    logic [7:0] sub_a, sub_b;
    logic [8:0] sub_result;
    sequence sub_sequence;
        (flash_data == {8'h61, sub_a}) ##DELAY
        (flash_data == {8'h62, sub_b}) ##DELAY
        (flash_data == 16'h9312);// SUM
    endsequence

    logic [7:0] sub_a_reg, sub_b_reg;
    bus_shift #(.DELAY(5), .WIDTH(8)) sub_a_shifting (
        .clk(clk),
        .arst_n(arst_n),
        .in(sub_a),
        .out(sub_a_reg)
    );
    bus_shift #(.DELAY(3), .WIDTH(8)) sub_b_shifting (
        .clk(clk),
        .arst_n(arst_n),
        .in(sub_b),
        .out(sub_b_reg)
    );

    assign sub_result = sub_a_reg - sub_b_reg;

    property p_exec_sub_from_reset;
    @(posedge clk) disable iff (!arst_n)
        $rose(arst_n) |-> sub_sequence |=> (alu_opcode==3'b001 && alu_result==sub_result[7:0]);
    endproperty


    // =============================== JMP assert BlackBox 
    logic [11:0] next_jump, next_jump_reg;
    bus_shift #(.DELAY(3), .WIDTH(12)) next_jump_shifting (
        .clk(clk),
        .arst_n(arst_n),
        .in(next_jump),
        .out(next_jump_reg)
    );

    sequence jmp_sequence;
        (flash_data == {4'h3, next_jump}) ##DELAY // JMP
        (flash_data == 16'h0000); // NOP
    endsequence

    property p_exec_jmp_from_reset;
    @(posedge clk) disable iff (!arst_n)
        $rose(arst_n) |->  jmp_sequence |=> (pc_out == next_jump_reg);
    endproperty


    // =============================== BC assert BlackBox 
    logic [7:0] carry_a, carry_b;
    sequence bc_sequence;
        (flash_data == {8'h61, carry_a}) ##DELAY
        (flash_data == {8'h62, carry_b}) ##DELAY
        (flash_data == 16'h8312) ##DELAY // SUM
        (flash_data == {4'h5, next_jump}) ##DELAY // BC
        (flash_data == 16'h0000);
    endsequence

    logic [7:0] carry_a_reg, carry_b_reg;
    bus_shift #(.DELAY(9), .WIDTH(8)) carry_a_shifting (
        .clk(clk),
        .arst_n(arst_n),
        .in(carry_a),
        .out(carry_a_reg)
    );
    bus_shift #(.DELAY(7), .WIDTH(8)) carry_b_shifting (
        .clk(clk),
        .arst_n(arst_n),
        .in(carry_b),
        .out(carry_b_reg)
    );

    logic [8:0] carry_result;
    assign carry_result = carry_b_reg + carry_a_reg;

    assume property (@(posedge clk) disable iff (!arst_n)
        bc_sequence |=> carry_result[8]);

    property p_exec_branch_carry_from_reset;
    @(posedge clk) disable iff (!arst_n)
        $rose(arst_n) |-> bc_sequence |=> (carry_result[8] && pc_out==next_jump_reg);
    endproperty

    // =============================== BEQ assert BlackBox 
    logic [7:0] cmp_a, cmp_b;
    sequence beq_sequence;
        (flash_data == {8'h61, cmp_a}) ##DELAY
        (flash_data == {8'h62, cmp_b}) ##DELAY
        (flash_data == 16'hD012) ##DELAY // CMP
        (flash_data == {4'h4, next_jump})  ##DELAY // BEQ
        (flash_data == 16'h0000); 
    endsequence

    logic [7:0] cmp_a_reg, cmp_b_reg;
    bus_shift #(.DELAY(9), .WIDTH(8)) cmp_a_shifting (
        .clk(clk),
        .arst_n(arst_n),
        .in(cmp_a),
        .out(cmp_a_reg)
    );
    bus_shift #(.DELAY(7), .WIDTH(8)) cmp_b_shifting (
        .clk(clk),
        .arst_n(arst_n),
        .in(cmp_b),
        .out(cmp_b_reg)
    );

    assume property (@(posedge clk) disable iff (!arst_n)
        1'b1 |-> cmp_a_reg == cmp_b_reg);

    property p_exec_branch_equal_from_reset;
    @(posedge clk) disable iff (!arst_n)
        $rose(arst_n) |-> beq_sequence |=> (pc_out==next_jump_reg);
    endproperty


    // =============================== IN-STORE assert BlackBox 

    sequence in_sequence;
        (flash_data == 16'h3200) ##DELAY
        (flash_data == 16'h6100) ##DELAY
        (flash_data == 16'h2101);// SUM
    endsequence

    logic [7:0] in_reg;
    bus_shift #(.DELAY(3), .WIDTH(8)) in_shifting (
        .clk(clk),
        .arst_n(arst_n),
        .in(in),
        .out(in_reg)
    ); 

    assume property (@(posedge clk) disable iff (!arst_n)
    1'b1 |-> cmp_a_reg == cmp_b_reg);

    property p_exec_in_from_reset;
    @(posedge clk) disable iff (!arst_n)
        $rose(arst_n) |-> in_sequence |=> sram_addr == 1'b1 |-> (in_reg == sram_data_in);
    endproperty

    // ============================ WhiteBox: suma y carry
    logic [8:0] sum;
    logic msb_sum_reg;
    assign sum = alu_a + alu_b;

    `AST(ALU, add,
        (alu_opcode == 3'b000) |->,
        (alu_result == sum[7:0] && carry_out == sum[8])
    )

    shift #(DELAY) carry_shifthing (
        .clk(clk),
        .arst_n(arst_n),
        .in(sum[8]),
        .out(msb_sum_reg)
    );

    `AST(ALU, carry_out,
        (alu_opcode == 3'b000) |-> ##DELAY,
        (carry_flag == msb_sum_reg)
    )

uC_ast_ADD:   assert property (p_exec_sum_from_reset);
uC_ast_SUB:   assert property (p_exec_sub_from_reset);
uC_ast_JMP:   assert property (p_exec_jmp_from_reset);
uC_ast_BC:    assert property (p_exec_branch_carry_from_reset);
uC_ast_BEQ:   assert property (p_exec_branch_equal_from_reset);
uC_ast_IN:    assert property (p_exec_in_from_reset);


endmodule

bind uC_8bits fv_uC_8bits fv_uC_8bits_i(.*);
